`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:49:54 12/31/2024 
// Design Name: 
// Module Name:    instructionMem 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module instructionMem(PC,out);

input [7:0] PC;
output reg [15:0] out;
 
reg [15:0] ROM [255:0];

initial 
begin

	ROM [0]  = 16'b001001_000_000_0110;		// li $t0,9					// 9
   ROM [1]  = 16'b000010_000_001_0110;		// li $t1,2					// 2
   ROM [2]  = 16'b000_001_000_010_0000;	// add $t2,$t0,$t1		// 11
	ROM [3] = 16'b001010_000_010_0101;		// addi $t2,$t0,10   	// 19
   ROM [4]  = 16'b010_000_000_010_0001;	// sll $t2,$t0,$t1		// 36
   ROM [5]  = 16'b010_000_000_010_0010;	// srl $t2,$t0,$t1		// 2
   ROM [6]  = 16'b000_001_000_010_1101;	// mul $t2,$t0,$t1		// 18
   ROM [7]  = 16'b000_001_000_010_0011;	// or $t2,$t0,$t1			// 11
   ROM [8]  = 16'b000_001_000_010_0100;	// and $t2,$t0,$t1		// 0
	
   ROM [9]  = 16'b110010_000_011_0110;		// li $t3,50				// 50
   ROM [10]  = 16'b000_011_011_100_1101;	// mul $t4,$t3,$t3		// 2500
   ROM [11] = 16'b000_100_011_101_1101;	// mul $t5,$t4,$t3		// 59464
	
   ROM [12] = 16'b000000_000_010_1100;		// mflo $t2					// 1
   ROM [13] = 16'b000000_000_010_1110;		// mfhi $t2					// 59464

	ROM [14] = 16'b001001_000_000_0110;		// li $t0,9
	ROM [15] = 16'b001010_000_010_0110;		// li $t2,10
	ROM [16] = 16'b000000_000_001_0110;		// li $t1,0
														// loop:
	ROM [17] = 16'b000001_001_001_0101; 	// addi $t1,$t1,1
	ROM [18] = 16'b000_001_000_011_1101;	// mul $t3,$t0,$t1
	ROM [19] = 16'b000000_001_011_1000;		// sw $t3,0($t1)
	ROM [20] = 16'b011000_010_001_1011;		// beq $t1,$t2,exit
														
	ROM [21] = 16'b000_000010001_1001;		// j loop
	
	ROM [22] = 16'b001001_000_000_0110;
	ROM [23] = 16'b001001_000_000_0110;
   ROM [24] = 16'b001001_000_000_0110;
														// exit:
	ROM [25] = 16'b000001_000_000_0110;		// li $t0,1
	ROM [26] = 16'b001010_000_010_0110;		// li $t2,10
	
														// loop2:
	ROM [27] = 16'b000000_010_001_0111;		// lw $t1,0($t2)
	ROM [28] = 16'b100001_000_010_1011;		// beq $t2,$t0,exit2
	ROM [29] = 16'b000_000_010_010_1111;	// sub $t2,$t2,$t0
	ROM [30] = 16'b000_000011011_1001;		// j loop2
	 
	ROM [31] = 16'b001001_000_000_0110;		
	ROM [32] = 16'b001001_000_000_0110;	
														// exit2:
														// rest all li $t0,9
	ROM [33] = 16'b001001_000_000_0110;
   ROM [34] = 16'b001001_000_000_0110;
   ROM [35] = 16'b001001_000_000_0110;
   ROM [36] = 16'b001001_000_000_0110;
   ROM [37] = 16'b001001_000_000_0110;
   ROM [38] = 16'b001001_000_000_0110;
   ROM [39] = 16'b001001_000_000_0110;
   ROM [40] = 16'b001001_000_000_0110;
   ROM [41] = 16'b001001_000_000_0110;
   ROM [42] = 16'b001001_000_000_0110;
   ROM [43] = 16'b001001_000_000_0110;
   ROM [44] = 16'b001001_000_000_0110;
   ROM [45] = 16'b001001_000_000_0110;
   ROM [46] = 16'b001001_000_000_0110;
   ROM [47] = 16'b001001_000_000_0110;
   ROM [48] = 16'b001001_000_000_0110;
   ROM [49] = 16'b001001_000_000_0110;
   ROM [50] = 16'b001001_000_000_0110;
   ROM [51] = 16'b001001_000_000_0110;
   ROM [52] = 16'b001001_000_000_0110;
   ROM [53] = 16'b001001_000_000_0110;
   ROM [54] = 16'b001001_000_000_0110;
   ROM [55] = 16'b001001_000_000_0110;
   ROM [56] = 16'b001001_000_000_0110;
   ROM [57] = 16'b001001_000_000_0110;
   ROM [58] = 16'b001001_000_000_0110;
   ROM [59] = 16'b001001_000_000_0110;
   ROM [60] = 16'b001001_000_000_0110;
   ROM [61] = 16'b001001_000_000_0110;
   ROM [62] = 16'b001001_000_000_0110;
   ROM [63] = 16'b001001_000_000_0110;
   ROM [64] = 16'b001001_000_000_0110;
   ROM [65] = 16'b001001_000_000_0110;
   ROM [66] = 16'b001001_000_000_0110;
   ROM [67] = 16'b001001_000_000_0110;
   ROM [68] = 16'b001001_000_000_0110;
   ROM [69] = 16'b001001_000_000_0110;
   ROM [70] = 16'b001001_000_000_0110;
   ROM [71] = 16'b001001_000_000_0110;
   ROM [72] = 16'b001001_000_000_0110;
   ROM [73] = 16'b001001_000_000_0110;
   ROM [74] = 16'b001001_000_000_0110;
   ROM [75] = 16'b001001_000_000_0110;
   ROM [76] = 16'b001001_000_000_0110;
   ROM [77] = 16'b001001_000_000_0110;
   ROM [78] = 16'b001001_000_000_0110;
   ROM [79] = 16'b001001_000_000_0110;
   ROM [80] = 16'b001001_000_000_0110;
   ROM [81] = 16'b001001_000_000_0110;
   ROM [82] = 16'b001001_000_000_0110;
   ROM [83] = 16'b001001_000_000_0110;
   ROM [84] = 16'b001001_000_000_0110;
   ROM [85] = 16'b001001_000_000_0110;
   ROM [86] = 16'b001001_000_000_0110;
   ROM [87] = 16'b001001_000_000_0110;
   ROM [88] = 16'b001001_000_000_0110;
   ROM [89] = 16'b001001_000_000_0110;
   ROM [90] = 16'b001001_000_000_0110;
   ROM [91] = 16'b001001_000_000_0110;
   ROM [92] = 16'b001001_000_000_0110;
   ROM [93] = 16'b001001_000_000_0110;
   ROM [94] = 16'b001001_000_000_0110;
   ROM [95] = 16'b001001_000_000_0110;
   ROM [96] = 16'b001001_000_000_0110;
   ROM [97] = 16'b001001_000_000_0110;
   ROM [98] = 16'b001001_000_000_0110;
   ROM [99] = 16'b001001_000_000_0110;
   ROM [100] = 16'b001001_000_000_0110;
   ROM [101] = 16'b001001_000_000_0110;
   ROM [102] = 16'b001001_000_000_0110;
   ROM [103] = 16'b001001_000_000_0110;
   ROM [104] = 16'b001001_000_000_0110;
   ROM [105] = 16'b001001_000_000_0110;
   ROM [106] = 16'b001001_000_000_0110;
   ROM [107] = 16'b001001_000_000_0110;
   ROM [108] = 16'b001001_000_000_0110;
   ROM [109] = 16'b001001_000_000_0110;
   ROM [110] = 16'b001001_000_000_0110;
   ROM [111] = 16'b001001_000_000_0110;
   ROM [112] = 16'b001001_000_000_0110;
   ROM [113] = 16'b001001_000_000_0110;
   ROM [114] = 16'b001001_000_000_0110;
   ROM [115] = 16'b001001_000_000_0110;
   ROM [116] = 16'b001001_000_000_0110;
   ROM [117] = 16'b001001_000_000_0110;
   ROM [118] = 16'b001001_000_000_0110;
   ROM [119] = 16'b001001_000_000_0110;
   ROM [120] = 16'b001001_000_000_0110;
   ROM [121] = 16'b001001_000_000_0110;
   ROM [122] = 16'b001001_000_000_0110;
   ROM [123] = 16'b001001_000_000_0110;
   ROM [124] = 16'b001001_000_000_0110;
   ROM [125] = 16'b001001_000_000_0110;
   ROM [126] = 16'b001001_000_000_0110;
   ROM [127] = 16'b001001_000_000_0110;
   ROM [128] = 16'b001001_000_000_0110;
   ROM [129] = 16'b001001_000_000_0110;
   ROM [130] = 16'b001001_000_000_0110;
   ROM [131] = 16'b001001_000_000_0110;
   ROM [132] = 16'b001001_000_000_0110;
   ROM [133] = 16'b001001_000_000_0110;
   ROM [134] = 16'b001001_000_000_0110;
   ROM [135] = 16'b001001_000_000_0110;
   ROM [136] = 16'b001001_000_000_0110;
   ROM [137] = 16'b001001_000_000_0110;
   ROM [138] = 16'b001001_000_000_0110;
   ROM [139] = 16'b001001_000_000_0110;
   ROM [140] = 16'b001001_000_000_0110;
   ROM [141] = 16'b001001_000_000_0110;
   ROM [142] = 16'b001001_000_000_0110;
   ROM [143] = 16'b001001_000_000_0110;
   ROM [144] = 16'b001001_000_000_0110;
   ROM [145] = 16'b001001_000_000_0110;
   ROM [146] = 16'b001001_000_000_0110;
   ROM [147] = 16'b001001_000_000_0110;
   ROM [148] = 16'b001001_000_000_0110;
   ROM [149] = 16'b001001_000_000_0110;
   ROM [150] = 16'b001001_000_000_0110;
   ROM [151] = 16'b001001_000_000_0110;
   ROM [152] = 16'b001001_000_000_0110;
   ROM [153] = 16'b001001_000_000_0110;
   ROM [154] = 16'b001001_000_000_0110;
   ROM [155] = 16'b001001_000_000_0110;
   ROM [156] = 16'b001001_000_000_0110;
   ROM [157] = 16'b001001_000_000_0110;
   ROM [158] = 16'b001001_000_000_0110;
   ROM [159] = 16'b001001_000_000_0110;
   ROM [160] = 16'b001001_000_000_0110;
   ROM [161] = 16'b001001_000_000_0110;
   ROM [162] = 16'b001001_000_000_0110;
   ROM [163] = 16'b001001_000_000_0110;
   ROM [164] = 16'b001001_000_000_0110;
   ROM [165] = 16'b001001_000_000_0110;
   ROM [166] = 16'b001001_000_000_0110;
   ROM [167] = 16'b001001_000_000_0110;
   ROM [168] = 16'b001001_000_000_0110;
   ROM [169] = 16'b001001_000_000_0110;
   ROM [170] = 16'b001001_000_000_0110;
   ROM [171] = 16'b001001_000_000_0110;
   ROM [172] = 16'b001001_000_000_0110;
   ROM [173] = 16'b001001_000_000_0110;
   ROM [174] = 16'b001001_000_000_0110;
   ROM [175] = 16'b001001_000_000_0110;
   ROM [176] = 16'b001001_000_000_0110;
   ROM [177] = 16'b001001_000_000_0110;
   ROM [178] = 16'b001001_000_000_0110;
   ROM [179] = 16'b001001_000_000_0110;
   ROM [180] = 16'b001001_000_000_0110;
   ROM [181] = 16'b001001_000_000_0110;
   ROM [182] = 16'b001001_000_000_0110;
   ROM [183] = 16'b001001_000_000_0110;
   ROM [184] = 16'b001001_000_000_0110;
   ROM [185] = 16'b001001_000_000_0110;
   ROM [186] = 16'b001001_000_000_0110;
   ROM [187] = 16'b001001_000_000_0110;
   ROM [188] = 16'b001001_000_000_0110;
   ROM [189] = 16'b001001_000_000_0110;
   ROM [190] = 16'b001001_000_000_0110;
   ROM [191] = 16'b001001_000_000_0110;
   ROM [192] = 16'b001001_000_000_0110;
   ROM [193] = 16'b001001_000_000_0110;
   ROM [194] = 16'b001001_000_000_0110;
   ROM [195] = 16'b001001_000_000_0110;
   ROM [196] = 16'b001001_000_000_0110;
   ROM [197] = 16'b001001_000_000_0110;
   ROM [198] = 16'b001001_000_000_0110;
   ROM [199] = 16'b001001_000_000_0110;
   ROM [200] = 16'b001001_000_000_0110;
   ROM [201] = 16'b001001_000_000_0110;
   ROM [202] = 16'b001001_000_000_0110;
   ROM [203] = 16'b001001_000_000_0110;
   ROM [204] = 16'b001001_000_000_0110;
   ROM [205] = 16'b001001_000_000_0110;
   ROM [206] = 16'b001001_000_000_0110;
   ROM [207] = 16'b001001_000_000_0110;
   ROM [208] = 16'b001001_000_000_0110;
   ROM [209] = 16'b001001_000_000_0110;
   ROM [210] = 16'b001001_000_000_0110;
   ROM [211] = 16'b001001_000_000_0110;
   ROM [212] = 16'b001001_000_000_0110;
   ROM [213] = 16'b001001_000_000_0110;
   ROM [214] = 16'b001001_000_000_0110;
   ROM [215] = 16'b001001_000_000_0110;
   ROM [216] = 16'b001001_000_000_0110;
   ROM [217] = 16'b001001_000_000_0110;
   ROM [218] = 16'b001001_000_000_0110;
   ROM [219] = 16'b001001_000_000_0110;
   ROM [220] = 16'b001001_000_000_0110;
   ROM [221] = 16'b001001_000_000_0110;
   ROM [222] = 16'b001001_000_000_0110;
   ROM [223] = 16'b001001_000_000_0110;
   ROM [224] = 16'b001001_000_000_0110;
   ROM [225] = 16'b001001_000_000_0110;
   ROM [226] = 16'b001001_000_000_0110;
   ROM [227] = 16'b001001_000_000_0110;
   ROM [228] = 16'b001001_000_000_0110;
   ROM [229] = 16'b001001_000_000_0110;
   ROM [230] = 16'b001001_000_000_0110;
   ROM [231] = 16'b001001_000_000_0110;
   ROM [232] = 16'b001001_000_000_0110;
   ROM [233] = 16'b001001_000_000_0110;
   ROM [234] = 16'b001001_000_000_0110;
   ROM [235] = 16'b001001_000_000_0110;
   ROM [236] = 16'b001001_000_000_0110;
   ROM [237] = 16'b001001_000_000_0110;
   ROM [238] = 16'b001001_000_000_0110;
   ROM [239] = 16'b001001_000_000_0110;
   ROM [240] = 16'b001001_000_000_0110;
   ROM [241] = 16'b001001_000_000_0110;
   ROM [242] = 16'b001001_000_000_0110;
   ROM [243] = 16'b001001_000_000_0110;
   ROM [244] = 16'b001001_000_000_0110;
   ROM [245] = 16'b001001_000_000_0110;
   ROM [246] = 16'b001001_000_000_0110;
   ROM [247] = 16'b001001_000_000_0110;
   ROM [248] = 16'b001001_000_000_0110;
   ROM [249] = 16'b001001_000_000_0110;
   ROM [250] = 16'b001001_000_000_0110;
   ROM [251] = 16'b001001_000_000_0110;
   ROM [252] = 16'b001001_000_000_0110;
   ROM [253] = 16'b001001_000_000_0110;
   ROM [254] = 16'b001001_000_000_0110;
   ROM [255] = 16'b001001_000_000_0110;

end

always @ (PC)
begin
	out = ROM[PC];
end

endmodule
